library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

use work.Lan9254Pkg.all;
use work.Lan9254ESCPkg.all;

entity Lan9254ESCrun is
end entity Lan9254ESCrun;

architecture rtl of Lan9254ESCrun is
   signal clk      : std_logic := '0';
   signal rst      : std_logic := '0';
   signal run      : boolean   := true;

   signal req      : Lan9254ReqType := LAN9254REQ_INIT_C;
   signal rep      : Lan9254RepType := LAN9254REP_INIT_C;

   signal al       : std_logic_vector(31 downto 0) := x"0000_0002";
   signal as       : std_logic_vector(31 downto 0) := x"0000_0001";

   signal cnt      : integer := 0;

   signal rxPDOMst : Lan9254PDOMstType;
   signal rxPDORdy : std_logic;

   signal txPDOMst : Lan9254PDOMstType := LAN9254PDO_MST_INIT_C;
   signal txPDORdy : std_logic;

begin

   process is begin
      if ( run ) then
         wait for 10 us;
         clk <= not clk;
      else
         wait;
      end if;
   end process;

   txPDOMst.ben   <= "11";

   process ( clk ) is
   begin
      if ( rising_edge( clk ) ) then
         if ( txPDOMst.valid = '0' ) then
            txPDOMst.data    <= (others => '0');
            txPDOMst.wrdAddr <= (others => '0');
            txPDOMst.valid   <= '1';
         elsif ( txPDORdy = '1' ) then
            txPDOMst.data    <= std_logic_vector(to_unsigned(cnt, txPDOMst.data'length));
            cnt              <= cnt + 1;
            txPDOMst.wrdAddr <= txPDOMst.wrdAddr + 1;
            if ( txPDOMst.wrdAddr >= unsigned(ESC_SM3_LEN_C) ) then
               txPDOMst.wrdAddr <= (others => '0');
            end if;
         end if;
      end if;
   end process;

   U_DUT : entity work.Lan9254ESC
      port map (
         clk         => clk,
         rst         => rst,

         req         => req,
         rep         => rep,

         rxPdoMst    => rxPDOMst,
         rxPdoRdy    => rxPDORdy,

         txPDOMst    => txPDOMst,
         txPDORdy    => txPDORdy
      );

   U_HBI : entity work.Lan9254Hbi
      generic map (
         CLOCK_FREQ_G => 12.0E6
      )
      port map (
         clk         => clk,
         rst         => rst,
         req         => req,
         rep         => rep
      );

   U_RXPDO : entity work.RxPDOSoft
      port map (
         clk         => clk,
         rst         => rst,

         rxPdoMst    => rxPDOMst,
         rxPdoRdy    => rxPDORdy

      );

end architecture rtl;
